VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR3B
  CLASS BLOCK ;
  FOREIGN NOR3B ;
  ORIGIN 0.770 0.420 ;
  SIZE 9.630 BY 3.040 ;
  OBS
      LAYER nwell ;
        RECT 6.930 2.200 8.860 2.380 ;
        RECT -0.180 -0.180 2.700 1.990 ;
      LAYER pwell ;
        RECT 3.200 -0.180 3.840 1.890 ;
      LAYER nwell ;
        RECT 4.740 1.210 8.860 2.200 ;
        RECT 6.910 0.760 8.860 1.210 ;
      LAYER pwell ;
        RECT 4.790 -0.130 6.880 0.550 ;
        RECT 7.240 -0.180 8.860 0.600 ;
      LAYER li1 ;
        RECT -0.770 0.900 -0.290 1.230 ;
        RECT 0.000 1.100 2.520 2.600 ;
        RECT 2.930 1.870 4.500 2.040 ;
        RECT 2.930 1.200 3.100 1.870 ;
        RECT 3.330 1.400 3.990 1.700 ;
        RECT 2.930 0.900 3.650 1.200 ;
        RECT -0.770 0.170 -0.290 0.500 ;
        RECT 2.930 0.300 3.100 0.900 ;
        RECT 3.820 0.650 3.990 1.400 ;
        RECT 4.330 1.050 4.500 1.870 ;
        RECT 4.920 1.390 5.630 2.600 ;
        RECT 5.880 1.220 6.180 2.020 ;
        RECT 6.430 1.390 6.730 2.600 ;
        RECT 5.880 1.050 6.730 1.220 ;
        RECT 4.330 0.720 5.350 1.050 ;
        RECT 0.000 0.000 3.100 0.300 ;
        RECT 3.280 -0.400 3.990 0.650 ;
        RECT 6.130 0.550 6.380 0.880 ;
        RECT 6.560 0.850 6.730 1.050 ;
        RECT 7.410 0.940 8.120 2.600 ;
        RECT 6.560 0.520 7.240 0.850 ;
        RECT 4.980 -0.400 5.630 0.420 ;
        RECT 6.560 0.380 6.730 0.520 ;
        RECT 6.430 0.000 6.730 0.380 ;
        RECT 7.470 -0.400 8.120 0.420 ;
        RECT 8.370 0.000 8.670 2.200 ;
      LAYER met1 ;
        RECT -0.180 2.220 8.850 2.620 ;
        RECT 0.000 -0.420 8.850 -0.020 ;
  END
END NOR3B
END LIBRARY

