magic
tech sky130A
timestamp 1757784183
<< nwell >>
rect 695 224 840 225
rect -79 81 3464 224
rect 1042 80 1315 81
rect 1455 80 1615 81
rect 2346 80 2591 81
rect 2782 80 3355 81
<< nmos >>
rect 0 0 15 42
rect 300 0 315 42
rect 600 -40 615 2
rect 960 -40 975 2
rect 1300 0 1315 42
rect 1600 0 1615 42
rect 1900 0 1915 42
rect 2260 -40 2275 2
rect 2700 -40 2715 2
rect 3040 0 3055 42
rect 3340 0 3355 42
<< pmos >>
rect 0 100 15 205
rect 300 100 315 205
rect 600 100 615 205
rect 960 100 975 205
rect 1300 100 1315 205
rect 1600 100 1615 205
rect 1900 100 1915 205
rect 2260 100 2275 205
rect 2700 100 2715 205
rect 3040 100 3055 205
rect 3340 100 3355 205
<< ndiff >>
rect -60 30 0 42
rect -60 12 -42 30
rect -20 12 0 30
rect -60 0 0 12
rect 15 30 75 42
rect 15 12 35 30
rect 57 12 75 30
rect 15 0 75 12
rect 240 30 300 42
rect 240 12 258 30
rect 280 12 300 30
rect 240 0 300 12
rect 315 30 375 42
rect 315 12 335 30
rect 357 12 375 30
rect 315 0 375 12
rect 540 -10 600 2
rect 540 -28 558 -10
rect 580 -28 600 -10
rect 540 -40 600 -28
rect 615 -10 675 2
rect 615 -28 635 -10
rect 657 -28 675 -10
rect 615 -40 675 -28
rect 1240 30 1300 42
rect 1240 12 1258 30
rect 1280 12 1300 30
rect 900 -10 960 2
rect 900 -28 918 -10
rect 940 -28 960 -10
rect 900 -40 960 -28
rect 975 -10 1035 2
rect 1240 0 1300 12
rect 1315 30 1375 42
rect 1315 12 1335 30
rect 1357 12 1375 30
rect 1315 0 1375 12
rect 1540 30 1600 42
rect 1540 12 1558 30
rect 1580 12 1600 30
rect 1540 0 1600 12
rect 1615 30 1675 42
rect 1615 12 1635 30
rect 1657 12 1675 30
rect 1615 0 1675 12
rect 1840 30 1900 42
rect 1840 12 1858 30
rect 1880 12 1900 30
rect 1840 0 1900 12
rect 1915 30 1975 42
rect 1915 12 1935 30
rect 1957 12 1975 30
rect 1915 0 1975 12
rect 975 -28 995 -10
rect 1017 -28 1035 -10
rect 975 -40 1035 -28
rect 2200 -10 2260 2
rect 2200 -28 2218 -10
rect 2240 -28 2260 -10
rect 2200 -40 2260 -28
rect 2275 -10 2335 2
rect 2275 -28 2295 -10
rect 2317 -28 2335 -10
rect 2275 -40 2335 -28
rect 2980 30 3040 42
rect 2980 12 2998 30
rect 3020 12 3040 30
rect 2640 -10 2700 2
rect 2640 -28 2658 -10
rect 2680 -28 2700 -10
rect 2640 -40 2700 -28
rect 2715 -10 2775 2
rect 2980 0 3040 12
rect 3055 30 3115 42
rect 3055 12 3075 30
rect 3097 12 3115 30
rect 3055 0 3115 12
rect 3280 30 3340 42
rect 3280 12 3298 30
rect 3320 12 3340 30
rect 3280 0 3340 12
rect 3355 30 3415 42
rect 3355 12 3375 30
rect 3397 12 3415 30
rect 3355 0 3415 12
rect 2715 -28 2735 -10
rect 2757 -28 2775 -10
rect 2715 -40 2775 -28
<< pdiff >>
rect -60 191 0 205
rect -60 112 -42 191
rect -20 112 0 191
rect -60 100 0 112
rect 15 191 75 205
rect 15 112 34 191
rect 56 112 75 191
rect 15 100 75 112
rect 240 191 300 205
rect 240 112 258 191
rect 280 112 300 191
rect 240 100 300 112
rect 315 191 375 205
rect 315 112 334 191
rect 356 112 375 191
rect 540 191 600 205
rect 315 100 375 112
rect 540 112 558 191
rect 580 112 600 191
rect 540 100 600 112
rect 615 191 675 205
rect 615 112 634 191
rect 656 112 675 191
rect 900 191 960 205
rect 615 100 675 112
rect 900 112 918 191
rect 940 112 960 191
rect 900 100 960 112
rect 975 191 1035 205
rect 975 112 994 191
rect 1016 112 1035 191
rect 975 100 1035 112
rect 1240 191 1300 205
rect 1240 112 1258 191
rect 1280 112 1300 191
rect 1240 100 1300 112
rect 1315 191 1375 205
rect 1315 112 1334 191
rect 1356 112 1375 191
rect 1315 100 1375 112
rect 1540 191 1600 205
rect 1540 112 1558 191
rect 1580 112 1600 191
rect 1540 100 1600 112
rect 1615 191 1675 205
rect 1615 112 1634 191
rect 1656 112 1675 191
rect 1615 100 1675 112
rect 1840 191 1900 205
rect 1840 112 1858 191
rect 1880 112 1900 191
rect 1840 100 1900 112
rect 1915 191 1975 205
rect 1915 112 1934 191
rect 1956 112 1975 191
rect 2200 191 2260 205
rect 1915 100 1975 112
rect 2200 112 2218 191
rect 2240 112 2260 191
rect 2200 100 2260 112
rect 2275 191 2335 205
rect 2275 112 2294 191
rect 2316 112 2335 191
rect 2640 191 2700 205
rect 2275 100 2335 112
rect 2640 112 2658 191
rect 2680 112 2700 191
rect 2640 100 2700 112
rect 2715 191 2775 205
rect 2715 112 2734 191
rect 2756 112 2775 191
rect 2715 100 2775 112
rect 2980 191 3040 205
rect 2980 112 2998 191
rect 3020 112 3040 191
rect 2980 100 3040 112
rect 3055 191 3115 205
rect 3055 112 3074 191
rect 3096 112 3115 191
rect 3055 100 3115 112
rect 3280 191 3340 205
rect 3280 112 3298 191
rect 3320 112 3340 191
rect 3280 100 3340 112
rect 3355 191 3415 205
rect 3355 112 3374 191
rect 3396 112 3415 191
rect 3355 100 3415 112
<< ndiffc >>
rect -42 12 -20 30
rect 35 12 57 30
rect 258 12 280 30
rect 335 12 357 30
rect 558 -28 580 -10
rect 635 -28 657 -10
rect 1258 12 1280 30
rect 918 -28 940 -10
rect 1335 12 1357 30
rect 1558 12 1580 30
rect 1635 12 1657 30
rect 1858 12 1880 30
rect 1935 12 1957 30
rect 995 -28 1017 -10
rect 2218 -28 2240 -10
rect 2295 -28 2317 -10
rect 2998 12 3020 30
rect 2658 -28 2680 -10
rect 3075 12 3097 30
rect 3298 12 3320 30
rect 3375 12 3397 30
rect 2735 -28 2757 -10
<< pdiffc >>
rect -42 112 -20 191
rect 34 112 56 191
rect 258 112 280 191
rect 334 112 356 191
rect 558 112 580 191
rect 634 112 656 191
rect 918 112 940 191
rect 994 112 1016 191
rect 1258 112 1280 191
rect 1334 112 1356 191
rect 1558 112 1580 191
rect 1634 112 1656 191
rect 1858 112 1880 191
rect 1934 112 1956 191
rect 2218 112 2240 191
rect 2294 112 2316 191
rect 2658 112 2680 191
rect 2734 112 2756 191
rect 2998 112 3020 191
rect 3074 112 3096 191
rect 3298 112 3320 191
rect 3374 112 3396 191
<< poly >>
rect 0 205 15 218
rect 300 205 315 218
rect 600 205 615 218
rect 960 205 975 218
rect 1300 205 1315 218
rect 1600 205 1615 218
rect 1900 205 1915 218
rect 2260 205 2275 218
rect 2700 205 2715 218
rect 3040 205 3055 218
rect 3340 205 3355 218
rect 473 145 515 153
rect 473 120 482 145
rect 505 120 515 145
rect 473 113 515 120
rect -129 77 -86 83
rect -129 49 -121 77
rect -95 71 -86 77
rect 0 71 15 100
rect -95 56 15 71
rect -95 49 -86 56
rect -129 43 -86 49
rect 0 42 15 56
rect 171 77 214 83
rect 171 49 179 77
rect 205 71 214 77
rect 300 71 315 100
rect 482 92 502 113
rect 826 145 871 153
rect 826 119 835 145
rect 861 119 871 145
rect 826 110 871 119
rect 600 92 615 100
rect 482 76 615 92
rect 832 88 861 110
rect 2122 142 2162 149
rect 2122 120 2130 142
rect 2153 120 2162 142
rect 2122 114 2162 120
rect 960 88 975 100
rect 832 73 975 88
rect 1171 77 1214 83
rect 832 72 961 73
rect 205 56 315 71
rect 205 49 214 56
rect 171 43 214 49
rect 300 42 315 56
rect 1171 49 1179 77
rect 1205 71 1214 77
rect 1300 71 1315 100
rect 1205 56 1315 71
rect 1205 49 1214 56
rect 1171 43 1214 49
rect 1300 42 1315 56
rect 1471 77 1514 83
rect 1471 49 1479 77
rect 1505 71 1514 77
rect 1600 71 1615 100
rect 1505 56 1615 71
rect 1505 49 1514 56
rect 1471 43 1514 49
rect 1600 42 1615 56
rect 1771 77 1814 83
rect 1771 49 1779 77
rect 1805 71 1814 77
rect 1900 71 1915 100
rect 1805 56 1915 71
rect 2131 85 2152 114
rect 2566 145 2611 153
rect 2566 119 2575 145
rect 2601 119 2611 145
rect 2566 110 2611 119
rect 2260 85 2275 100
rect 2131 69 2275 85
rect 2572 88 2601 110
rect 2700 88 2715 100
rect 2572 73 2715 88
rect 2911 77 2954 83
rect 2572 72 2701 73
rect 1805 49 1814 56
rect 1771 43 1814 49
rect 1900 42 1915 56
rect 2911 49 2919 77
rect 2945 71 2954 77
rect 3040 71 3055 100
rect 2945 56 3055 71
rect 2945 49 2954 56
rect 2911 43 2954 49
rect 3040 42 3055 56
rect 3211 77 3254 83
rect 3211 49 3219 77
rect 3245 71 3254 77
rect 3340 71 3355 100
rect 3245 56 3355 71
rect 3245 49 3254 56
rect 3211 43 3254 49
rect 3340 42 3355 56
rect 502 15 615 34
rect 0 -13 15 0
rect 300 -13 315 0
rect 502 -2 527 15
rect 600 2 615 15
rect 818 14 975 31
rect 818 8 837 14
rect 470 -10 527 -2
rect 470 -27 478 -10
rect 495 -27 527 -10
rect 470 -34 527 -27
rect 470 -35 502 -34
rect 794 0 837 8
rect 960 2 975 14
rect 794 -28 802 0
rect 830 -28 837 0
rect 794 -36 837 -28
rect 2136 11 2275 26
rect 2136 3 2154 11
rect 1300 -13 1315 0
rect 1600 -13 1615 0
rect 1900 -13 1915 0
rect 2109 -6 2154 3
rect 2260 2 2275 11
rect 2558 14 2715 31
rect 2558 8 2577 14
rect 2109 -32 2118 -6
rect 2145 -32 2154 -6
rect 2109 -40 2154 -32
rect 2534 0 2577 8
rect 2700 2 2715 14
rect 2534 -28 2542 0
rect 2570 -28 2577 0
rect 2534 -36 2577 -28
rect 3040 -13 3055 0
rect 3340 -13 3355 0
rect 600 -53 615 -40
rect 960 -53 975 -40
rect 2260 -53 2275 -40
rect 2700 -53 2715 -40
<< polycont >>
rect 482 120 505 145
rect -121 49 -95 77
rect 179 49 205 77
rect 835 119 861 145
rect 2130 120 2153 142
rect 1179 49 1205 77
rect 1479 49 1505 77
rect 1779 49 1805 77
rect 2575 119 2601 145
rect 2919 49 2945 77
rect 3219 49 3245 77
rect 478 -27 495 -10
rect 802 -28 830 0
rect 2118 -32 2145 -6
rect 2542 -28 2570 0
<< locali >>
rect -143 246 92 249
rect -143 226 -42 246
rect -19 226 92 246
rect 162 246 392 249
rect 162 226 258 246
rect 281 226 392 246
rect 464 246 692 249
rect 464 226 558 246
rect 581 226 692 246
rect 824 246 1052 249
rect 824 226 918 246
rect 941 226 1052 246
rect 1162 246 1392 249
rect 1162 226 1258 246
rect 1281 226 1392 246
rect 1462 246 1692 249
rect 1462 226 1558 246
rect 1581 226 1692 246
rect 1762 246 1992 249
rect 1762 226 1858 246
rect 1881 226 1992 246
rect 2124 246 2352 249
rect 2124 226 2218 246
rect 2241 226 2352 246
rect 2564 246 2792 249
rect 2564 226 2658 246
rect 2681 226 2792 246
rect 2902 246 3132 249
rect 2902 226 2998 246
rect 3021 226 3132 246
rect 3202 246 3432 249
rect 3202 226 3298 246
rect 3321 226 3432 246
rect -49 199 -13 226
rect 251 199 287 226
rect 1251 199 1287 226
rect 1551 199 1587 226
rect 1851 199 1887 226
rect 2991 199 3027 226
rect 3291 199 3327 226
rect -50 191 -11 199
rect -143 143 -99 147
rect -143 121 -132 143
rect -108 121 -99 143
rect -143 118 -99 121
rect -50 112 -42 191
rect -20 112 -11 191
rect -50 106 -11 112
rect 25 191 64 199
rect 25 112 34 191
rect 56 112 64 191
rect 250 191 289 199
rect 126 141 151 146
rect 126 120 130 141
rect 147 120 151 141
rect 126 119 151 120
rect 25 106 64 112
rect -129 77 -86 83
rect -129 76 -121 77
rect -143 51 -121 76
rect -129 49 -121 51
rect -95 49 -86 77
rect -129 43 -86 49
rect 33 73 55 106
rect 127 76 149 119
rect 250 112 258 191
rect 280 112 289 191
rect 250 106 289 112
rect 325 191 364 199
rect 325 112 334 191
rect 356 112 364 191
rect 550 191 589 199
rect 473 145 515 153
rect 473 140 482 145
rect 325 106 364 112
rect 430 120 482 140
rect 505 120 515 145
rect 430 118 515 120
rect 171 77 214 83
rect 171 76 179 77
rect 72 73 94 75
rect 33 56 75 73
rect 92 56 94 73
rect 33 36 55 56
rect 72 53 94 56
rect 127 51 179 76
rect 171 49 179 51
rect 205 49 214 77
rect 171 43 214 49
rect 333 73 355 106
rect 381 94 413 96
rect 381 73 385 94
rect 333 68 385 73
rect 411 73 413 94
rect 430 73 452 118
rect 473 113 515 118
rect 550 112 558 191
rect 580 112 589 191
rect 550 106 589 112
rect 625 191 664 199
rect 625 112 634 191
rect 656 112 664 191
rect 910 191 949 199
rect 826 146 871 153
rect 727 145 871 146
rect 727 143 835 145
rect 727 121 733 143
rect 756 121 835 143
rect 727 119 835 121
rect 861 119 871 145
rect 727 117 871 119
rect 625 106 664 112
rect 826 110 871 117
rect 910 112 918 191
rect 940 112 949 191
rect 910 106 949 112
rect 985 191 1024 199
rect 985 112 994 191
rect 1016 112 1024 191
rect 985 106 1024 112
rect 1250 191 1289 199
rect 1250 112 1258 191
rect 1280 112 1289 191
rect 1250 106 1289 112
rect 1325 191 1364 199
rect 1325 112 1334 191
rect 1356 112 1364 191
rect 1325 106 1364 112
rect 1550 191 1589 199
rect 1550 112 1558 191
rect 1580 112 1589 191
rect 1550 106 1589 112
rect 1625 191 1664 199
rect 1625 112 1634 191
rect 1656 112 1664 191
rect 1850 191 1889 199
rect 1625 106 1664 112
rect 1722 142 1763 145
rect 1722 106 1726 142
rect 1759 106 1763 142
rect 1850 112 1858 191
rect 1880 112 1889 191
rect 1850 106 1889 112
rect 1925 191 1964 199
rect 1925 112 1934 191
rect 1956 112 1964 191
rect 2093 193 2122 197
rect 2093 170 2097 193
rect 2118 176 2156 193
rect 2118 170 2122 176
rect 2093 166 2122 170
rect 2139 149 2156 176
rect 2210 191 2249 199
rect 2122 142 2162 149
rect 2122 120 2130 142
rect 2153 120 2162 142
rect 2122 114 2162 120
rect 1925 106 1964 112
rect 2210 112 2218 191
rect 2240 112 2249 191
rect 2210 106 2249 112
rect 2285 191 2324 199
rect 2285 112 2294 191
rect 2316 112 2324 191
rect 2650 191 2689 199
rect 2566 145 2611 153
rect 2285 106 2324 112
rect 2420 139 2454 142
rect 2420 112 2424 139
rect 2450 138 2454 139
rect 2566 138 2575 145
rect 2450 119 2575 138
rect 2601 119 2611 145
rect 2450 118 2611 119
rect 2450 112 2454 118
rect 2420 108 2454 112
rect 2566 110 2611 118
rect 2650 112 2658 191
rect 2680 112 2689 191
rect 2650 106 2689 112
rect 2725 191 2764 199
rect 2725 112 2734 191
rect 2756 112 2764 191
rect 2725 106 2764 112
rect 2990 191 3029 199
rect 2990 112 2998 191
rect 3020 112 3029 191
rect 2990 106 3029 112
rect 3065 191 3104 199
rect 3065 112 3074 191
rect 3096 112 3104 191
rect 3065 106 3104 112
rect 3290 191 3329 199
rect 3290 112 3298 191
rect 3320 112 3329 191
rect 3290 106 3329 112
rect 3365 191 3404 199
rect 3365 112 3374 191
rect 3396 112 3404 191
rect 3365 106 3404 112
rect 411 68 451 73
rect 333 56 451 68
rect 333 36 355 56
rect 556 51 583 106
rect -52 30 -9 36
rect -52 12 -42 30
rect -20 12 -9 30
rect -52 6 -9 12
rect 24 30 67 36
rect 24 12 35 30
rect 57 12 67 30
rect 24 6 67 12
rect 248 30 291 36
rect 248 12 258 30
rect 280 12 291 30
rect 248 6 291 12
rect 324 30 367 36
rect 324 12 335 30
rect 357 12 367 30
rect 387 35 411 39
rect 387 18 391 35
rect 408 34 411 35
rect 468 34 583 51
rect 408 18 485 34
rect 387 16 485 18
rect 324 6 367 12
rect -45 -17 -21 6
rect 255 -17 279 6
rect 420 -7 451 -5
rect -142 -19 83 -17
rect -142 -36 -44 -19
rect -23 -36 83 -19
rect -142 -40 83 -36
rect 165 -19 383 -17
rect 165 -36 256 -19
rect 277 -36 383 -19
rect 420 -25 428 -7
rect 446 -12 451 -7
rect 470 -10 502 -2
rect 556 -4 583 34
rect 633 73 655 106
rect 633 69 786 73
rect 633 56 751 69
rect 633 -4 655 56
rect 746 36 751 56
rect 780 36 786 69
rect 746 32 786 36
rect 916 30 943 106
rect 710 9 746 14
rect 470 -12 478 -10
rect 446 -25 478 -12
rect 420 -27 478 -25
rect 495 -27 502 -10
rect 420 -29 502 -27
rect 470 -35 502 -29
rect 548 -10 591 -4
rect 548 -28 558 -10
rect 580 -28 591 -10
rect 548 -34 591 -28
rect 624 -10 667 -4
rect 624 -28 635 -10
rect 657 -28 667 -10
rect 710 -18 716 9
rect 740 1 746 9
rect 857 13 943 30
rect 794 1 837 8
rect 740 0 837 1
rect 740 -18 802 0
rect 710 -19 802 -18
rect 710 -22 746 -19
rect 624 -34 667 -28
rect 794 -28 802 -19
rect 830 -28 837 0
rect 794 -36 837 -28
rect 165 -40 383 -36
rect 857 -56 876 13
rect 916 -4 943 13
rect 993 73 1015 106
rect 1171 77 1214 83
rect 993 63 1059 73
rect 1096 67 1127 70
rect 1171 67 1179 77
rect 1096 66 1179 67
rect 1096 63 1100 66
rect 993 56 1100 63
rect 993 -4 1015 56
rect 1042 46 1100 56
rect 1096 42 1100 46
rect 1122 49 1179 66
rect 1205 49 1214 77
rect 1122 42 1127 49
rect 1171 43 1214 49
rect 1333 73 1355 106
rect 1397 78 1431 81
rect 1397 73 1401 78
rect 1333 56 1401 73
rect 1096 39 1127 42
rect 1333 36 1355 56
rect 1397 51 1401 56
rect 1427 73 1431 78
rect 1471 77 1514 83
rect 1471 73 1479 77
rect 1427 56 1479 73
rect 1427 51 1431 56
rect 1397 48 1431 51
rect 1471 49 1479 56
rect 1505 49 1514 77
rect 1471 43 1514 49
rect 1633 73 1655 106
rect 1722 102 1763 106
rect 1727 100 1758 102
rect 1683 74 1706 77
rect 1683 73 1686 74
rect 1633 56 1686 73
rect 1703 56 1706 74
rect 1633 36 1655 56
rect 1683 53 1706 56
rect 1727 76 1754 100
rect 1771 77 1814 83
rect 1771 76 1779 77
rect 1727 51 1779 76
rect 1771 49 1779 51
rect 1805 49 1814 77
rect 1771 43 1814 49
rect 1933 73 1955 106
rect 1933 59 2079 73
rect 2216 59 2243 106
rect 1933 56 2243 59
rect 1933 36 1955 56
rect 2062 42 2243 56
rect 1248 30 1291 36
rect 1248 12 1258 30
rect 1280 12 1291 30
rect 1248 6 1291 12
rect 1324 30 1367 36
rect 1324 12 1335 30
rect 1357 12 1367 30
rect 1324 6 1367 12
rect 1548 30 1591 36
rect 1548 12 1558 30
rect 1580 12 1591 30
rect 1548 6 1591 12
rect 1624 30 1667 36
rect 1624 12 1635 30
rect 1657 12 1667 30
rect 1624 6 1667 12
rect 1848 30 1891 36
rect 1848 12 1858 30
rect 1880 12 1891 30
rect 1848 6 1891 12
rect 1924 30 1967 36
rect 1924 12 1935 30
rect 1957 12 1967 30
rect 1924 6 1967 12
rect 908 -10 951 -4
rect 908 -28 918 -10
rect 940 -28 951 -10
rect 908 -34 951 -28
rect 984 -10 1027 -4
rect 984 -28 995 -10
rect 1017 -28 1027 -10
rect 984 -34 1027 -28
rect 849 -60 878 -56
rect 849 -78 854 -60
rect 873 -78 878 -60
rect 849 -82 878 -78
rect 1255 -107 1279 6
rect 1555 -107 1579 6
rect 1855 -107 1879 6
rect 2109 -6 2154 3
rect 2216 -4 2243 42
rect 2293 73 2315 106
rect 2293 69 2526 73
rect 2293 56 2491 69
rect 2293 -4 2315 56
rect 2486 36 2491 56
rect 2520 36 2526 69
rect 2486 32 2526 36
rect 2656 30 2683 106
rect 2597 13 2683 30
rect 2356 1 2387 5
rect 2534 1 2577 8
rect 2109 -21 2118 -6
rect 2065 -25 2118 -21
rect 2015 -29 2118 -25
rect 2015 -56 2019 -29
rect 2048 -32 2118 -29
rect 2145 -32 2154 -6
rect 2048 -38 2154 -32
rect 2208 -10 2251 -4
rect 2208 -28 2218 -10
rect 2240 -28 2251 -10
rect 2208 -34 2251 -28
rect 2284 -10 2327 -4
rect 2284 -28 2295 -10
rect 2317 -28 2327 -10
rect 2356 -20 2361 1
rect 2382 0 2577 1
rect 2382 -19 2542 0
rect 2382 -20 2387 -19
rect 2356 -24 2387 -20
rect 2284 -34 2327 -28
rect 2534 -28 2542 -19
rect 2570 -28 2577 0
rect 2534 -36 2577 -28
rect 2048 -44 2082 -38
rect 2109 -40 2154 -38
rect 2048 -56 2053 -44
rect 2597 -56 2616 13
rect 2656 -4 2683 13
rect 2733 73 2755 106
rect 2911 77 2954 83
rect 2733 63 2799 73
rect 2836 67 2867 70
rect 2911 67 2919 77
rect 2836 66 2919 67
rect 2836 63 2840 66
rect 2733 56 2840 63
rect 2733 -4 2755 56
rect 2782 46 2840 56
rect 2836 42 2840 46
rect 2862 49 2919 66
rect 2945 49 2954 77
rect 2862 42 2867 49
rect 2911 43 2954 49
rect 3073 73 3095 106
rect 3211 77 3254 83
rect 3211 73 3219 77
rect 3073 56 3219 73
rect 2836 39 2867 42
rect 3073 36 3095 56
rect 3211 49 3219 56
rect 3245 49 3254 77
rect 3211 43 3254 49
rect 3373 73 3395 106
rect 3423 74 3446 77
rect 3423 73 3426 74
rect 3373 56 3426 73
rect 3443 56 3464 74
rect 3373 36 3395 56
rect 3423 53 3446 56
rect 2988 30 3031 36
rect 2988 12 2998 30
rect 3020 12 3031 30
rect 2988 6 3031 12
rect 3064 30 3107 36
rect 3064 12 3075 30
rect 3097 12 3107 30
rect 3064 6 3107 12
rect 3288 30 3331 36
rect 3288 12 3298 30
rect 3320 12 3331 30
rect 3288 6 3331 12
rect 3364 30 3407 36
rect 3364 12 3375 30
rect 3397 12 3407 30
rect 3364 6 3407 12
rect 2648 -10 2691 -4
rect 2648 -28 2658 -10
rect 2680 -28 2691 -10
rect 2648 -34 2691 -28
rect 2724 -10 2767 -4
rect 2724 -28 2735 -10
rect 2757 -28 2767 -10
rect 2724 -34 2767 -28
rect 2015 -60 2053 -56
rect 2589 -60 2618 -56
rect 2589 -78 2594 -60
rect 2613 -78 2618 -60
rect 2589 -82 2618 -78
rect 2995 -107 3019 6
rect 3295 -107 3319 6
rect 465 -109 683 -107
rect 465 -126 556 -109
rect 577 -126 683 -109
rect 465 -130 683 -126
rect 825 -109 1043 -107
rect 825 -126 916 -109
rect 937 -126 1043 -109
rect 825 -130 1043 -126
rect 1165 -109 1383 -107
rect 1165 -126 1256 -109
rect 1277 -126 1383 -109
rect 1165 -130 1383 -126
rect 1465 -109 1683 -107
rect 1465 -126 1556 -109
rect 1577 -126 1683 -109
rect 1465 -130 1683 -126
rect 1765 -109 1983 -107
rect 1765 -126 1856 -109
rect 1877 -126 1983 -109
rect 1765 -130 1983 -126
rect 2125 -109 2343 -107
rect 2125 -126 2216 -109
rect 2237 -126 2343 -109
rect 2125 -130 2343 -126
rect 2565 -109 2783 -107
rect 2565 -126 2656 -109
rect 2677 -126 2783 -109
rect 2565 -130 2783 -126
rect 2905 -109 3123 -107
rect 2905 -126 2996 -109
rect 3017 -126 3123 -109
rect 2905 -130 3123 -126
rect 3205 -109 3423 -107
rect 3205 -126 3296 -109
rect 3317 -126 3423 -109
rect 3205 -130 3423 -126
<< viali >>
rect -42 226 -19 246
rect 258 226 281 246
rect 558 226 581 246
rect 918 226 941 246
rect 1258 226 1281 246
rect 1558 226 1581 246
rect 1858 226 1881 246
rect 2218 226 2241 246
rect 2658 226 2681 246
rect 2998 226 3021 246
rect 3298 226 3321 246
rect -132 121 -108 143
rect 130 120 147 141
rect 75 56 92 73
rect 385 68 411 94
rect 733 121 756 143
rect 1726 106 1759 142
rect 2097 170 2118 193
rect 2424 112 2450 139
rect 391 18 408 35
rect -44 -36 -23 -19
rect 256 -36 277 -19
rect 428 -25 446 -7
rect 751 36 780 69
rect 716 -18 740 9
rect 1100 42 1122 66
rect 1401 51 1427 78
rect 1686 56 1703 74
rect 854 -78 873 -60
rect 2491 36 2520 69
rect 2019 -56 2048 -29
rect 2361 -20 2382 1
rect 2840 42 2862 66
rect 3426 56 3443 74
rect 2594 -78 2613 -60
rect 556 -126 577 -109
rect 916 -126 937 -109
rect 1256 -126 1277 -109
rect 1556 -126 1577 -109
rect 1856 -126 1877 -109
rect 2216 -126 2237 -109
rect 2656 -126 2677 -109
rect 2996 -126 3017 -109
rect 3296 -126 3317 -109
<< metal1 >>
rect -143 246 3464 255
rect -143 226 -42 246
rect -19 226 258 246
rect 281 226 558 246
rect 581 226 918 246
rect 941 226 1258 246
rect 1281 226 1558 246
rect 1581 226 1858 246
rect 1881 226 2218 246
rect 2241 226 2658 246
rect 2681 226 2998 246
rect 3021 226 3298 246
rect 3321 226 3464 246
rect -143 220 3464 226
rect 1991 219 2139 220
rect 2335 219 2455 220
rect 2089 193 2125 200
rect 2089 191 2097 193
rect 727 171 2097 191
rect 727 152 765 171
rect 2089 170 2097 171
rect 2118 191 2125 193
rect 2118 171 2373 191
rect 2118 170 2125 171
rect 2089 163 2125 170
rect -143 143 765 152
rect -143 121 -132 143
rect -108 141 733 143
rect -108 121 130 141
rect -143 120 130 121
rect 147 121 733 141
rect 756 121 765 143
rect 147 120 765 121
rect -143 113 765 120
rect 1719 142 1765 147
rect 379 94 417 98
rect 65 77 95 80
rect 65 73 112 77
rect 65 56 75 73
rect 92 56 112 73
rect 379 68 385 94
rect 411 68 417 94
rect 379 64 417 68
rect 65 49 112 56
rect 95 37 112 49
rect 387 37 414 41
rect 95 35 414 37
rect 95 18 391 35
rect 408 18 414 35
rect 95 13 414 18
rect 387 12 414 13
rect 434 -2 456 113
rect 1719 106 1726 142
rect 1759 106 1765 142
rect 1719 100 1765 106
rect 1394 78 1434 84
rect 742 69 791 78
rect 742 36 751 69
rect 780 67 791 69
rect 1090 67 1134 74
rect 780 66 1134 67
rect 780 42 1100 66
rect 1122 42 1134 66
rect 1394 51 1401 78
rect 1427 51 1434 78
rect 1394 45 1434 51
rect 1678 74 1709 82
rect 1678 56 1686 74
rect 1703 56 1709 74
rect 1678 48 1709 56
rect 780 37 1134 42
rect 780 36 791 37
rect 742 28 791 36
rect 416 -7 456 -2
rect -142 -19 398 -9
rect -142 -36 -44 -19
rect -23 -36 256 -19
rect 277 -36 398 -19
rect 416 -25 428 -7
rect 446 -25 456 -7
rect 710 9 746 14
rect 710 -18 716 9
rect 742 -18 746 9
rect 710 -22 746 -18
rect 1688 -20 1705 48
rect 416 -32 456 -25
rect -142 -44 398 -36
rect 362 -99 398 -44
rect 1101 -34 1705 -20
rect 2353 8 2373 171
rect 2416 139 2458 145
rect 2416 112 2424 139
rect 2450 112 2458 139
rect 2416 105 2458 112
rect 2482 69 2531 78
rect 3418 74 3449 82
rect 2482 36 2491 69
rect 2520 67 2531 69
rect 2830 67 2874 74
rect 2520 66 2874 67
rect 2520 42 2840 66
rect 2862 42 2874 66
rect 3418 56 3426 74
rect 3443 56 3449 74
rect 3418 48 3449 56
rect 2520 37 2874 42
rect 2520 36 2531 37
rect 2482 28 2531 36
rect 2353 1 2389 8
rect 2353 -20 2361 1
rect 2382 -20 2389 1
rect 3428 -20 3445 48
rect 2009 -29 2058 -22
rect 2353 -27 2389 -20
rect 845 -60 882 -53
rect 845 -78 854 -60
rect 873 -66 882 -60
rect 1101 -66 1118 -34
rect 2009 -56 2019 -29
rect 2048 -56 2058 -29
rect 2841 -34 3445 -20
rect 2009 -64 2058 -56
rect 2585 -60 2622 -53
rect 873 -78 1118 -66
rect 845 -80 1118 -78
rect 2585 -78 2594 -60
rect 2613 -66 2622 -60
rect 2841 -66 2858 -34
rect 2613 -78 2858 -66
rect 2585 -80 2858 -78
rect 845 -85 882 -80
rect 2585 -85 2622 -80
rect 2353 -99 2501 -98
rect 362 -109 3459 -99
rect 362 -126 556 -109
rect 577 -126 916 -109
rect 937 -126 1256 -109
rect 1277 -126 1556 -109
rect 1577 -126 1856 -109
rect 1877 -126 2216 -109
rect 2237 -126 2656 -109
rect 2677 -126 2996 -109
rect 3017 -126 3296 -109
rect 3317 -126 3459 -109
rect 362 -134 3459 -126
<< via1 >>
rect 385 68 411 94
rect 1726 106 1759 142
rect 1401 51 1427 78
rect 716 -18 740 9
rect 740 -18 742 9
rect 2424 112 2450 139
rect 2019 -56 2048 -29
<< metal2 >>
rect 1719 142 1765 147
rect 1719 134 1726 142
rect 1401 107 1726 134
rect 379 94 417 98
rect 379 68 385 94
rect 411 69 417 94
rect 1401 84 1427 107
rect 1719 106 1726 107
rect 1759 106 1765 142
rect 1719 100 1765 106
rect 2416 139 2458 145
rect 2416 112 2424 139
rect 2450 112 2458 139
rect 2416 105 2458 112
rect 1394 78 1434 84
rect 411 68 710 69
rect 379 64 710 68
rect 402 55 710 64
rect 695 14 710 55
rect 1394 51 1401 78
rect 1427 51 1434 78
rect 1394 45 1434 51
rect 695 9 746 14
rect 695 -18 716 9
rect 742 -18 746 9
rect 695 -22 746 -18
rect 721 -81 741 -22
rect 2009 -29 2058 -22
rect 2009 -56 2019 -29
rect 2048 -56 2058 -29
rect 2009 -64 2058 -56
rect 2024 -81 2041 -64
rect 2416 -81 2436 105
rect 721 -95 2436 -81
<< labels >>
rlabel locali -143 62 -143 62 7 D
port 1 w
rlabel metal1 -143 237 -143 237 7 Vdd
port 3 w
rlabel metal1 -142 -30 -142 -30 7 GND
port 4 w
rlabel metal1 -143 132 -143 132 7 CLK
port 5 w
rlabel locali 3160 73 3160 73 1 Q
port 2 n
<< end >>
