magic
tech sky130A
timestamp 1756285088
<< nwell >>
rect -34 -18 117 149
<< pwell >>
rect -26 -104 109 -42
<< nmos >>
rect 34 -94 49 -52
<< pmos >>
rect 34 0 49 131
<< ndiff >>
rect -16 -63 34 -52
rect -16 -83 -7 -63
rect 10 -83 34 -63
rect -16 -94 34 -83
rect 49 -62 99 -52
rect 49 -82 76 -62
rect 93 -82 99 -62
rect 49 -94 99 -82
<< pdiff >>
rect -16 114 34 131
rect -16 13 -6 114
rect 11 13 34 114
rect -16 0 34 13
rect 49 110 99 131
rect 49 5 74 110
rect 91 5 99 110
rect 49 0 99 5
<< ndiffc >>
rect -7 -83 10 -63
rect 76 -82 93 -62
<< pdiffc >>
rect -6 13 11 114
rect 74 5 91 110
<< poly >>
rect 34 131 49 144
rect -69 -12 -35 -11
rect 34 -12 49 0
rect -69 -19 49 -12
rect -69 -36 -61 -19
rect -44 -36 49 -19
rect -69 -42 49 -36
rect -69 -43 -35 -42
rect 34 -52 49 -42
rect 34 -107 49 -94
<< polycont >>
rect -61 -36 -44 -19
<< locali >>
rect -15 163 20 171
rect -34 146 -20 163
rect -2 146 32 163
rect 50 146 92 163
rect 110 146 117 163
rect -15 114 20 146
rect -15 13 -6 114
rect 11 13 20 114
rect -15 5 20 13
rect 65 110 100 125
rect 65 5 74 110
rect 91 5 100 110
rect -69 -19 -35 -11
rect -69 -36 -61 -19
rect -44 -36 -35 -19
rect -69 -43 -35 -36
rect -15 -63 20 -55
rect -15 -83 -7 -63
rect 10 -83 20 -63
rect -15 -109 20 -83
rect 65 -62 100 5
rect 65 -82 76 -62
rect 93 -82 100 -62
rect 65 -91 100 -82
rect -25 -126 -17 -109
rect 0 -126 33 -109
rect 50 -126 89 -109
rect 106 -126 109 -109
<< viali >>
rect -20 146 -2 163
rect 32 146 50 163
rect 92 146 110 163
rect -17 -126 0 -109
rect 33 -126 50 -109
rect 89 -126 106 -109
<< metal1 >>
rect -34 163 117 173
rect -34 146 -20 163
rect -2 146 32 163
rect 50 146 92 163
rect 110 146 117 163
rect -34 133 117 146
rect -26 -109 109 -97
rect -26 -126 -17 -109
rect 0 -126 33 -109
rect 50 -126 89 -109
rect 106 -126 109 -109
rect -26 -137 109 -126
<< labels >>
rlabel polycont -61 -36 -44 -19 1 INPUT
rlabel locali 75 -37 92 -20 1 OUTPUT
rlabel metal1 60 -126 77 -109 1 GND
rlabel metal1 8 -126 25 -109 1 GND
rlabel metal1 6 146 23 163 1 VDD
rlabel metal1 63 146 80 163 1 VDD
<< end >>
