magic
tech sky130A
timestamp 1757776277
<< nwell >>
rect 693 220 885 238
rect -18 -18 270 199
rect 474 121 885 220
rect 691 76 885 121
<< pwell >>
rect 320 -18 384 189
rect 479 -13 688 55
rect 724 -18 885 60
<< nmos >>
rect 328 125 370 140
rect 328 70 370 85
rect 568 0 583 42
rect 623 0 638 42
rect 817 0 832 42
<< pmos >>
rect 568 139 583 202
rect 623 139 638 202
rect 0 90 252 105
rect 817 94 832 220
rect 0 35 252 50
<< ndiff >>
rect 328 164 370 175
rect 328 147 341 164
rect 362 147 370 164
rect 328 140 370 147
rect 328 114 370 125
rect 328 97 336 114
rect 357 97 370 114
rect 328 85 370 97
rect 328 63 370 70
rect 328 46 340 63
rect 357 46 370 63
rect 328 35 370 46
rect 533 33 568 42
rect 533 8 540 33
rect 557 8 568 33
rect 533 0 568 8
rect 583 0 623 42
rect 638 30 673 42
rect 638 8 649 30
rect 666 8 673 30
rect 638 0 673 8
rect 782 34 817 42
rect 782 8 789 34
rect 806 8 817 34
rect 782 0 817 8
rect 832 37 867 42
rect 832 8 843 37
rect 860 8 867 37
rect 832 0 867 8
<< pdiff >>
rect 782 210 817 220
rect 533 192 568 202
rect 533 149 540 192
rect 557 149 568 192
rect 0 135 252 140
rect 0 118 8 135
rect 235 118 252 135
rect 0 105 252 118
rect 533 139 568 149
rect 583 192 623 202
rect 583 149 594 192
rect 611 149 623 192
rect 583 139 623 149
rect 638 192 673 202
rect 638 149 649 192
rect 666 149 673 192
rect 638 139 673 149
rect 0 50 252 90
rect 782 104 789 210
rect 806 104 817 210
rect 782 94 817 104
rect 832 210 867 220
rect 832 105 843 210
rect 860 105 867 210
rect 832 94 867 105
rect 0 22 252 35
rect 0 5 8 22
rect 235 5 252 22
rect 0 0 252 5
<< ndiffc >>
rect 341 147 362 164
rect 336 97 357 114
rect 340 46 357 63
rect 540 8 557 33
rect 649 8 666 30
rect 789 8 806 34
rect 843 8 860 37
<< pdiffc >>
rect 540 149 557 192
rect 8 118 235 135
rect 594 149 611 192
rect 649 149 666 192
rect 789 104 806 210
rect 843 105 860 210
rect 8 5 235 22
<< psubdiff >>
rect 328 29 370 35
rect 328 12 340 29
rect 357 12 370 29
rect 328 0 370 12
rect 494 33 533 42
rect 494 8 506 33
rect 523 8 533 33
rect 494 0 533 8
rect 743 34 782 42
rect 743 8 755 34
rect 772 8 782 34
rect 743 0 782 8
<< nsubdiff >>
rect 741 210 782 220
rect 492 192 533 202
rect 0 169 252 181
rect 0 152 8 169
rect 235 152 252 169
rect 0 140 252 152
rect 492 149 504 192
rect 521 149 533 192
rect 492 139 533 149
rect 741 104 753 210
rect 770 104 782 210
rect 741 94 782 104
<< psubdiffcont >>
rect 340 12 357 29
rect 506 8 523 33
rect 755 8 772 34
<< nsubdiffcont >>
rect 8 152 235 169
rect 504 149 521 192
rect 753 104 770 210
<< poly >>
rect 817 220 832 233
rect 568 202 583 215
rect 623 202 638 217
rect -59 115 -26 123
rect -59 98 -54 115
rect -37 105 -26 115
rect 269 125 328 140
rect 370 125 383 140
rect 269 105 284 125
rect -37 98 0 105
rect -59 90 0 98
rect 252 90 284 105
rect 568 105 583 139
rect 502 97 583 105
rect 305 70 328 85
rect 370 70 383 85
rect 502 80 514 97
rect 531 80 583 97
rect 623 88 638 139
rect 502 72 583 80
rect 305 50 320 70
rect -59 42 0 50
rect -59 25 -54 42
rect -37 35 0 42
rect 252 35 320 50
rect 568 42 583 72
rect 609 80 642 88
rect 609 63 617 80
rect 634 63 642 80
rect 609 55 642 63
rect 691 77 728 85
rect 691 60 701 77
rect 718 76 728 77
rect 817 76 832 94
rect 718 60 832 76
rect 691 59 832 60
rect 623 42 638 55
rect 691 52 728 59
rect 817 42 832 59
rect -37 25 -26 35
rect -59 17 -26 25
rect 568 -13 583 0
rect 623 -13 638 0
rect 817 -13 832 0
<< polycont >>
rect -54 98 -37 115
rect 514 80 531 97
rect -54 25 -37 42
rect 617 63 634 80
rect 701 60 718 77
<< locali >>
rect 0 249 252 260
rect 0 232 2 249
rect 19 232 70 249
rect 87 232 148 249
rect 165 232 216 249
rect 233 232 252 249
rect 0 169 252 232
rect 492 249 563 260
rect 492 232 494 249
rect 511 232 544 249
rect 561 232 563 249
rect 0 152 8 169
rect 235 152 252 169
rect 0 135 252 152
rect -77 115 -29 123
rect -77 98 -54 115
rect -37 98 -29 115
rect 0 118 8 135
rect 235 118 252 135
rect 0 110 252 118
rect 293 187 450 204
rect 293 120 310 187
rect 333 164 399 170
rect 333 147 341 164
rect 362 147 399 164
rect 333 140 399 147
rect 293 114 365 120
rect -77 90 -29 98
rect 293 97 336 114
rect 357 97 365 114
rect 293 90 365 97
rect -77 42 -29 50
rect -77 25 -54 42
rect -37 25 -29 42
rect 293 30 310 90
rect 382 65 399 140
rect 433 105 450 187
rect 492 192 563 232
rect 643 251 673 260
rect 643 234 650 251
rect 667 234 673 251
rect 492 149 504 192
rect 521 149 540 192
rect 557 149 563 192
rect 492 139 563 149
rect 588 192 618 202
rect 588 149 594 192
rect 611 149 618 192
rect 588 122 618 149
rect 643 192 673 234
rect 643 149 649 192
rect 666 149 673 192
rect 643 139 673 149
rect 741 249 812 260
rect 741 248 793 249
rect 741 231 743 248
rect 760 232 793 248
rect 810 232 812 249
rect 760 231 812 232
rect 741 210 812 231
rect 588 105 673 122
rect 433 97 535 105
rect 433 80 514 97
rect 531 80 535 97
rect 433 72 535 80
rect 613 80 638 88
rect -77 17 -29 25
rect 0 22 310 30
rect 0 5 8 22
rect 235 5 310 22
rect 0 0 310 5
rect 328 63 399 65
rect 328 46 340 63
rect 357 46 399 63
rect 613 63 617 80
rect 634 63 638 80
rect 613 55 638 63
rect 656 85 673 105
rect 741 104 753 210
rect 770 104 789 210
rect 806 104 812 210
rect 741 94 812 104
rect 837 210 867 220
rect 837 105 843 210
rect 860 105 867 210
rect 656 77 724 85
rect 656 60 701 77
rect 718 60 724 77
rect 328 29 399 46
rect 656 52 724 60
rect 328 12 340 29
rect 357 12 399 29
rect 328 -12 399 12
rect 328 -29 330 -12
rect 347 -29 380 -12
rect 397 -29 399 -12
rect 328 -40 399 -29
rect 498 33 563 42
rect 656 38 673 52
rect 498 8 506 33
rect 523 8 540 33
rect 557 8 563 33
rect 498 -12 563 8
rect 643 30 673 38
rect 643 8 649 30
rect 666 8 673 30
rect 643 0 673 8
rect 747 34 812 42
rect 747 8 755 34
rect 772 8 789 34
rect 806 8 812 34
rect 498 -29 500 -12
rect 517 -29 544 -12
rect 561 -29 563 -12
rect 498 -40 563 -29
rect 747 -12 812 8
rect 837 37 867 105
rect 837 8 843 37
rect 860 8 867 37
rect 837 0 867 8
rect 747 -29 749 -12
rect 766 -29 793 -12
rect 810 -29 812 -12
rect 747 -40 812 -29
<< viali >>
rect 2 232 19 249
rect 70 232 87 249
rect 148 232 165 249
rect 216 232 233 249
rect 494 232 511 249
rect 544 232 561 249
rect 650 234 667 251
rect 743 231 760 248
rect 793 232 810 249
rect 330 -29 347 -12
rect 380 -29 397 -12
rect 500 -29 517 -12
rect 544 -29 561 -12
rect 749 -29 766 -12
rect 793 -29 810 -12
<< metal1 >>
rect -18 251 885 262
rect -18 249 650 251
rect -18 232 2 249
rect 19 232 70 249
rect 87 232 148 249
rect 165 232 216 249
rect 233 232 494 249
rect 511 232 544 249
rect 561 234 650 249
rect 667 249 885 251
rect 667 248 793 249
rect 667 234 743 248
rect 561 232 743 234
rect -18 231 743 232
rect 760 232 793 248
rect 810 232 885 249
rect 760 231 885 232
rect -18 222 885 231
rect 0 -12 885 -2
rect 0 -29 330 -12
rect 347 -29 380 -12
rect 397 -29 500 -12
rect 517 -29 544 -12
rect 561 -29 749 -12
rect 766 -29 793 -12
rect 810 -29 885 -12
rect 0 -42 885 -29
<< labels >>
rlabel metal1 428 -36 465 -8 1 gnd
rlabel metal1 666 -36 703 -8 1 gnd
rlabel metal1 72 -36 109 -8 1 gnd
rlabel metal1 -14 229 -4 253 1 vdd
rlabel metal1 344 232 384 257 1 vdd
rlabel metal1 576 226 616 251 1 vdd
rlabel metal1 839 231 879 256 1 vdd
rlabel locali 616 67 634 84 1 a
rlabel locali -74 98 -56 115 1 b
rlabel locali -73 25 -55 42 1 c
rlabel locali 844 58 862 75 1 out
rlabel locali 456 79 475 97 1 y0
rlabel locali 665 61 684 79 1 y1
rlabel pdiff 155 59 176 78 1 m
rlabel ndiff 593 10 614 29 1 n
<< end >>
