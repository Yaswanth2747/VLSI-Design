magic
tech sky130A
timestamp 1756296321
<< nwell >>
rect -22 225 62 239
rect -109 -77 111 225
<< pwell >>
rect -110 -268 112 -111
<< nmos >>
rect -14 -226 1 -142
<< pmos >>
rect -14 -57 1 205
<< ndiff >>
rect -47 -161 -14 -142
rect -47 -181 -39 -161
rect -22 -181 -14 -161
rect -47 -199 -14 -181
rect -47 -219 -39 -199
rect -22 -219 -14 -199
rect -47 -226 -14 -219
rect 1 -152 34 -142
rect 1 -172 9 -152
rect 26 -172 34 -152
rect 1 -190 34 -172
rect 1 -210 9 -190
rect 26 -210 34 -190
rect 1 -226 34 -210
<< pdiff >>
rect -47 165 -14 205
rect -47 145 -39 165
rect -22 145 -14 165
rect -47 93 -14 145
rect -47 73 -39 93
rect -22 73 -14 93
rect -47 5 -14 73
rect -47 -15 -39 5
rect -22 -15 -14 5
rect -47 -57 -14 -15
rect 1 179 34 205
rect 1 159 9 179
rect 26 159 34 179
rect 1 85 34 159
rect 1 65 9 85
rect 26 65 34 85
rect 1 -17 34 65
rect 1 -37 9 -17
rect 26 -37 34 -17
rect 1 -57 34 -37
<< ndiffc >>
rect -39 -181 -22 -161
rect -39 -219 -22 -199
rect 9 -172 26 -152
rect 9 -210 26 -190
<< pdiffc >>
rect -39 145 -22 165
rect -39 73 -22 93
rect -39 -15 -22 5
rect 9 159 26 179
rect 9 65 26 85
rect 9 -37 26 -17
<< poly >>
rect -14 205 1 218
rect -14 -86 1 -57
rect -144 -94 1 -86
rect -144 -112 -136 -94
rect -116 -112 1 -94
rect -144 -120 1 -112
rect -14 -142 1 -120
rect -14 -239 1 -226
<< polycont >>
rect -136 -112 -116 -94
<< locali >>
rect -49 225 -43 242
rect -26 225 -6 242
rect 11 225 45 242
rect -39 165 -22 225
rect -39 93 -22 145
rect -39 5 -22 73
rect -39 -49 -22 -15
rect 9 179 26 195
rect 9 85 26 159
rect 9 -17 26 65
rect -144 -94 -107 -86
rect -144 -112 -136 -94
rect -116 -112 -107 -94
rect -144 -120 -107 -112
rect -39 -161 -22 -151
rect -39 -199 -22 -181
rect 9 -152 26 -37
rect 9 -190 26 -172
rect 9 -218 26 -210
rect -39 -242 -22 -219
rect -54 -259 -39 -242
rect -22 -259 1 -242
rect 18 -259 40 -242
<< viali >>
rect -43 225 -26 242
rect -6 225 11 242
rect -39 -259 -22 -242
rect 1 -259 18 -242
<< metal1 >>
rect -54 242 53 246
rect -54 225 -43 242
rect -26 225 -6 242
rect 11 225 53 242
rect -54 214 53 225
rect -59 -242 48 -235
rect -59 -259 -39 -242
rect -22 -259 1 -242
rect 18 -259 48 -242
rect -59 -267 48 -259
<< labels >>
rlabel viali -43 225 -26 242 1 VDD
rlabel viali -6 225 11 242 1 VDD
rlabel viali -39 -259 -22 -242 1 GND
rlabel viali 1 -259 18 -242 1 GND
rlabel pdiffc 9 -37 26 -17 1 OUTPUT
rlabel pdiffc 9 65 26 85 1 OUTPUT
rlabel polycont -136 -112 -116 -94 1 INPUT
<< end >>
