* Assignment 1, Q2: INVX2 CMOS Inverter - DC VTC

.lib ~/VLSI_Design/open_pdks/sources/sky130_fd_pr/models/sky130.lib.spice tt

* parameters
.param VDD=1.8
.param Lmin=0.15
.param Wn1=0.42
.param Wp1=1.31   ; INVX1 widths
.param Wn2=0.84
.param Wp2=2.62   ; INVX2 widths = 2 * INVX1

.param ASn1=Wn1*0.3
.param ADn1=Wn1*0.3
.param PSn1=2*(Wn1+0.3)
.param PDn1=2*(Wn1+0.3)

.param ASp1=Wp1*0.3
.param ADp1=Wp1*0.3
.param PSp1=2*(Wp1+0.3)
.param PDp1=2*(Wp1+0.3)

.param ASn2=Wn2*0.3
.param ADn2=Wn2*0.3
.param PSn2=2*(Wn2+0.3)
.param PDn2=2*(Wn2+0.3)

.param ASp2=Wp2*0.3
.param ADp2=Wp2*0.3
.param PSp2=2*(Wp2+0.3)
.param PDp2=2*(Wp2+0.3)

Vdd vdd gnd DC {VDD}
Vin in gnd DC 0

* Main Circuit
Xinv2 in vdd gnd out INVX2_sub
Xload out vdd gnd out_load INVX1_sub

* Sub - Ckt Defn
.subckt INVX1_sub a vdd vss z
* NMOS
XM1 z a vss vss sky130_fd_pr__nfet_01v8 L={Lmin} W={Wn1} AS={ASn1} AD={ADn1} PS={PSn1} PD={PDn1}
* PMOS
XM2 z a vdd vdd sky130_fd_pr__pfet_01v8 L={Lmin} W={Wp1} AS={ASp1} AD={ADp1} PS={PSp1} PD={PDp1}
.ends INVX1_sub

.subckt INVX2_sub a vdd vss z
* NMOS
XM1 z a vss vss sky130_fd_pr__nfet_01v8 L={Lmin} W={Wn2} AS={ASn2} AD={ADn2} PS={PSn2} PD={PDn2}
* PMOS
XM2 z a vdd vdd sky130_fd_pr__pfet_01v8 L={Lmin} W={Wp2} AS={ASp2} AD={ADp2} PS={PSp2} PD={PDp2}
.ends INVX2_sub

.dc Vin 0 {VDD} 0.001

.control
run
set wr_singlescale
wrdata inverter_vtc_invx2.csv v(in) v(out)
plot v(out) vs v(in)
.endc

.end

