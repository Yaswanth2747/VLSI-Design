VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX1
  CLASS BLOCK ;
  FOREIGN INVX1 ;
  ORIGIN 0.910 1.360 ;
  SIZE 2.020 BY 3.040 ;
  OBS
      LAYER nwell ;
        RECT -0.600 -0.180 0.930 1.440 ;
      LAYER pwell ;
        RECT -0.180 -0.360 0.930 -0.340 ;
        RECT -0.480 -0.960 0.930 -0.360 ;
        RECT -0.180 -1.120 0.930 -0.960 ;
      LAYER li1 ;
        RECT -0.360 1.410 0.830 1.580 ;
        RECT -0.360 0.050 0.250 1.410 ;
        RECT 0.500 -0.160 0.750 1.210 ;
        RECT -0.910 -0.360 0.120 -0.160 ;
        RECT 0.500 -0.360 1.110 -0.160 ;
        RECT -0.360 -1.080 0.250 -0.570 ;
        RECT 0.500 -0.910 0.750 -0.360 ;
        RECT -0.360 -1.260 0.610 -1.080 ;
      LAYER met1 ;
        RECT -0.600 1.280 0.930 1.680 ;
        RECT -0.480 -1.360 0.930 -0.960 ;
  END
END INVX1
END LIBRARY

