* NGSPICE file created from INVX2.ext - technology: sky130A
.subckt INVX2 INPUT VDD GND OUTPUT
X0 OUTPUT INPUT VDD w_n109_n77# sky130_fd_pr__pfet_01v8 ad=0.8646 pd=5.9 as=0.8646 ps=5.9 w=2.62 l=0.15
X1 OUTPUT INPUT GND SUB sky130_fd_pr__nfet_01v8 ad=0.2772 pd=2.34 as=0.2772 ps=2.34 w=0.84 l=0.15
C0 OUTPUT INPUT 0.04562f
C1 GND VDD 0.02096f
C2 VDD INPUT 0.03366f
C3 GND INPUT 0.02558f
C4 OUTPUT w_n109_n77# 0.03361f
C5 VDD w_n109_n77# 0.05152f
C6 GND w_n109_n77# 0.00634f
C7 INPUT w_n109_n77# 0.07565f
C8 OUTPUT VDD 0.17359f
C9 OUTPUT GND 0.06593f
C10 GND SUB 0.19469f
C11 OUTPUT SUB 0.16834f
C12 VDD SUB 0.22411f
C13 INPUT SUB 0.34933f
C14 w_n109_n77# SUB 0.81139f
.ends
