* Transient analysis of INVX2 with PEX
.lib ~/VLSI_Design/open_pdks/sources/sky130_fd_pr/models/sky130.lib.spice tt

* --------------------------
* Parameters
* --------------------------
.param VDD=1.8
.param Vhalf={VDD/2}

* --------------------------
* Power supply and input
* --------------------------
Vdd vdd gnd DC {VDD}
Vin in gnd PULSE(0 {VDD} 0p 20p 20p 1n 2n)

* --------------------------
* Include extracted netlist (PEX)
* --------------------------
.include invx1_pex.spice
.include invx2_pex.spice

* --------------------------
* Instantiate inverter + load
* --------------------------
Xinv1 in vdd gnd out INVX2
Xload out vdd gnd out_load INVX1

* --------------------------
* Transient simulation
* --------------------------
.tran 1ps 10ns 0 10p

* --------------------------
* Measurements
* --------------------------
.meas tran tr   TRIG v(out) VAL='0.1*VDD' RISE=1 TARG v(out) VAL='0.9*VDD' RISE=1
.meas tran tf   TRIG v(out) VAL='0.9*VDD' FALL=1 TARG v(out) VAL='0.1*VDD' FALL=1
.meas tran tpHL TRIG v(in)  VAL='Vhalf'   RISE=1 TARG v(out) VAL='Vhalf' FALL=1
.meas tran tpLH TRIG v(in)  VAL='Vhalf'   FALL=1 TARG v(out) VAL='Vhalf' RISE=1

* --------------------------
* Control block
* --------------------------
.control
run
print tran tr tf tpHL tpLH
plot v(in) v(out)
.endc

.end

