* NGSPICE file created from INVX1.ext - technology: sky130A

.subckt INVX1 INPUT VDD GND OUTPUT
X0 OUTPUT INPUT GND SUB sky130_fd_pr__nfet_01v8 ad=0.21 pd=1.84 as=0.21 ps=1.84 w=0.42 l=0.15
**devattr s=2100,184 d=2100,184
X1 OUTPUT INPUT VDD w_n34_n18# sky130_fd_pr__pfet_01v8 ad=0.655 pd=3.62 as=0.655 ps=3.62 w=1.31 l=0.15
**devattr s=6550,362 d=6550,362
C0 w_n34_n18# GND 0.00611f
C1 VDD INPUT 0.03258f
C2 OUTPUT VDD 0.11449f
C3 OUTPUT INPUT 0.03339f
C4 GND VDD 0.04946f
C5 GND INPUT 0.02752f
C6 OUTPUT GND 0.07203f
C7 w_n34_n18# VDD 0.02841f
C8 w_n34_n18# INPUT 0.06021f
C9 OUTPUT w_n34_n18# 0.01037f
C10 GND SUB 0.21316f
C11 OUTPUT SUB 0.0978f
C12 VDD SUB 0.2575f
C13 INPUT SUB 0.27853f
C14 w_n34_n18# SUB 0.3026f
.ends

