VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dff
  CLASS BLOCK ;
  FOREIGN dff ;
  ORIGIN 1.430 1.340 ;
  SIZE 36.070 BY 3.890 ;
  PIN D
    ANTENNAGATEAREA 0.220500 ;
    PORT
      LAYER li1 ;
        RECT -1.290 0.760 -0.860 0.830 ;
        RECT -1.430 0.510 -0.860 0.760 ;
        RECT -1.290 0.430 -0.860 0.510 ;
    END
  END D
  PIN Q
    ANTENNAGATEAREA 0.220500 ;
    ANTENNADIFFAREA 0.882000 ;
    PORT
      LAYER li1 ;
        RECT 30.650 1.060 31.040 1.990 ;
        RECT 30.730 0.730 30.950 1.060 ;
        RECT 32.110 0.730 32.540 0.830 ;
        RECT 30.730 0.560 32.540 0.730 ;
        RECT 30.730 0.360 30.950 0.560 ;
        RECT 32.110 0.430 32.540 0.560 ;
        RECT 30.640 0.060 31.070 0.360 ;
    END
  END Q
  PIN Vdd
    ANTENNADIFFAREA 4.410000 ;
    PORT
      LAYER li1 ;
        RECT -1.430 2.260 0.920 2.490 ;
        RECT 1.620 2.260 3.920 2.490 ;
        RECT 4.640 2.260 6.920 2.490 ;
        RECT 8.240 2.260 10.520 2.490 ;
        RECT 11.620 2.260 13.920 2.490 ;
        RECT 14.620 2.260 16.920 2.490 ;
        RECT 17.620 2.260 19.920 2.490 ;
        RECT 21.240 2.260 23.520 2.490 ;
        RECT 25.640 2.260 27.920 2.490 ;
        RECT 29.020 2.260 31.320 2.490 ;
        RECT 32.020 2.260 34.320 2.490 ;
        RECT -0.490 1.990 -0.130 2.260 ;
        RECT 2.510 1.990 2.870 2.260 ;
        RECT 12.510 1.990 12.870 2.260 ;
        RECT 15.510 1.990 15.870 2.260 ;
        RECT 18.510 1.990 18.870 2.260 ;
        RECT 29.910 1.990 30.270 2.260 ;
        RECT 32.910 1.990 33.270 2.260 ;
        RECT -0.500 1.060 -0.110 1.990 ;
        RECT 2.500 1.060 2.890 1.990 ;
        RECT 12.500 1.060 12.890 1.990 ;
        RECT 15.500 1.060 15.890 1.990 ;
        RECT 18.500 1.060 18.890 1.990 ;
        RECT 29.900 1.060 30.290 1.990 ;
        RECT 32.900 1.060 33.290 1.990 ;
      LAYER met1 ;
        RECT -1.430 2.200 34.640 2.550 ;
        RECT 19.910 2.190 21.390 2.200 ;
        RECT 23.350 2.190 24.550 2.200 ;
    END
  END Vdd
  PIN GND
    ANTENNADIFFAREA 1.764000 ;
    PORT
      LAYER li1 ;
        RECT -0.520 0.060 -0.090 0.360 ;
        RECT 2.480 0.060 2.910 0.360 ;
        RECT 12.480 0.060 12.910 0.360 ;
        RECT 15.480 0.060 15.910 0.360 ;
        RECT 18.480 0.060 18.910 0.360 ;
        RECT 29.880 0.060 30.310 0.360 ;
        RECT 32.880 0.060 33.310 0.360 ;
        RECT -0.450 -0.170 -0.210 0.060 ;
        RECT 2.550 -0.170 2.790 0.060 ;
        RECT -1.420 -0.400 0.830 -0.170 ;
        RECT 1.650 -0.400 3.830 -0.170 ;
        RECT 12.550 -1.070 12.790 0.060 ;
        RECT 15.550 -1.070 15.790 0.060 ;
        RECT 18.550 -1.070 18.790 0.060 ;
        RECT 29.950 -1.070 30.190 0.060 ;
        RECT 32.950 -1.070 33.190 0.060 ;
        RECT 4.650 -1.300 6.830 -1.070 ;
        RECT 8.250 -1.300 10.430 -1.070 ;
        RECT 11.650 -1.300 13.830 -1.070 ;
        RECT 14.650 -1.300 16.830 -1.070 ;
        RECT 17.650 -1.300 19.830 -1.070 ;
        RECT 21.250 -1.300 23.430 -1.070 ;
        RECT 25.650 -1.300 27.830 -1.070 ;
        RECT 29.050 -1.300 31.230 -1.070 ;
        RECT 32.050 -1.300 34.230 -1.070 ;
      LAYER met1 ;
        RECT -1.420 -0.440 3.980 -0.090 ;
        RECT 3.620 -0.990 3.980 -0.440 ;
        RECT 23.530 -0.990 25.010 -0.980 ;
        RECT 3.620 -1.340 34.640 -0.990 ;
    END
  END GND
  PIN CLK
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 20.930 1.930 21.220 1.970 ;
        RECT 20.930 1.760 21.560 1.930 ;
        RECT 20.930 1.660 21.220 1.760 ;
        RECT -1.430 1.180 -0.990 1.470 ;
        RECT 8.260 1.460 8.710 1.530 ;
        RECT 21.390 1.490 21.560 1.760 ;
        RECT 1.260 1.190 1.510 1.460 ;
        RECT 1.270 0.760 1.490 1.190 ;
        RECT 7.270 1.170 8.710 1.460 ;
        RECT 8.260 1.100 8.710 1.170 ;
        RECT 21.220 1.140 21.620 1.490 ;
        RECT 1.710 0.760 2.140 0.830 ;
        RECT 1.270 0.510 2.140 0.760 ;
        RECT 1.710 0.430 2.140 0.510 ;
        RECT 23.560 0.010 23.870 0.050 ;
        RECT 25.340 0.010 25.770 0.080 ;
        RECT 4.200 -0.120 4.510 -0.050 ;
        RECT 4.700 -0.120 5.020 -0.020 ;
        RECT 4.200 -0.290 5.020 -0.120 ;
        RECT 23.560 -0.190 25.770 0.010 ;
        RECT 23.560 -0.240 23.870 -0.190 ;
        RECT 4.700 -0.350 5.020 -0.290 ;
        RECT 25.340 -0.360 25.770 -0.190 ;
      LAYER met1 ;
        RECT 20.890 1.910 21.250 2.000 ;
        RECT 7.270 1.710 23.730 1.910 ;
        RECT 7.270 1.520 7.650 1.710 ;
        RECT 20.890 1.630 21.250 1.710 ;
        RECT -1.430 1.130 7.650 1.520 ;
        RECT 4.340 -0.020 4.560 1.130 ;
        RECT 4.160 -0.320 4.560 -0.020 ;
        RECT 23.530 0.080 23.730 1.710 ;
        RECT 23.530 -0.270 23.890 0.080 ;
    END
  END CLK
  OBS
      LAYER nwell ;
        RECT 6.950 2.240 8.400 2.250 ;
        RECT -0.790 0.810 34.640 2.240 ;
        RECT 10.420 0.800 13.150 0.810 ;
        RECT 14.550 0.800 16.150 0.810 ;
        RECT 23.460 0.800 25.910 0.810 ;
        RECT 27.820 0.800 33.550 0.810 ;
      LAYER li1 ;
        RECT 0.250 1.060 0.640 1.990 ;
        RECT 3.250 1.060 3.640 1.990 ;
        RECT 4.730 1.400 5.150 1.530 ;
        RECT 4.300 1.180 5.150 1.400 ;
        RECT 0.330 0.730 0.550 1.060 ;
        RECT 0.720 0.730 0.940 0.750 ;
        RECT 0.330 0.560 0.940 0.730 ;
        RECT 0.330 0.360 0.550 0.560 ;
        RECT 0.720 0.530 0.940 0.560 ;
        RECT 3.330 0.730 3.550 1.060 ;
        RECT 3.810 0.730 4.130 0.960 ;
        RECT 4.300 0.730 4.520 1.180 ;
        RECT 4.730 1.130 5.150 1.180 ;
        RECT 5.500 1.060 5.890 1.990 ;
        RECT 6.250 1.060 6.640 1.990 ;
        RECT 9.100 1.060 9.490 1.990 ;
        RECT 9.850 1.060 10.240 1.990 ;
        RECT 13.250 1.060 13.640 1.990 ;
        RECT 16.250 1.060 16.640 1.990 ;
        RECT 3.330 0.560 4.510 0.730 ;
        RECT 3.330 0.360 3.550 0.560 ;
        RECT 5.560 0.510 5.830 1.060 ;
        RECT 0.240 0.060 0.670 0.360 ;
        RECT 3.240 0.060 3.670 0.360 ;
        RECT 3.870 0.340 4.110 0.390 ;
        RECT 4.680 0.340 5.830 0.510 ;
        RECT 3.870 0.160 4.850 0.340 ;
        RECT 5.560 -0.040 5.830 0.340 ;
        RECT 6.330 0.730 6.550 1.060 ;
        RECT 6.330 0.560 7.860 0.730 ;
        RECT 6.330 -0.040 6.550 0.560 ;
        RECT 7.460 0.320 7.860 0.560 ;
        RECT 9.160 0.300 9.430 1.060 ;
        RECT 7.100 0.010 7.460 0.140 ;
        RECT 8.570 0.130 9.430 0.300 ;
        RECT 7.940 0.010 8.370 0.080 ;
        RECT 5.480 -0.340 5.910 -0.040 ;
        RECT 6.240 -0.340 6.670 -0.040 ;
        RECT 7.100 -0.190 8.370 0.010 ;
        RECT 7.100 -0.220 7.460 -0.190 ;
        RECT 7.940 -0.360 8.370 -0.190 ;
        RECT 8.570 -0.560 8.760 0.130 ;
        RECT 9.160 -0.040 9.430 0.130 ;
        RECT 9.930 0.730 10.150 1.060 ;
        RECT 9.930 0.630 10.590 0.730 ;
        RECT 10.960 0.670 11.270 0.700 ;
        RECT 11.710 0.670 12.140 0.830 ;
        RECT 10.960 0.630 12.140 0.670 ;
        RECT 9.930 0.560 12.140 0.630 ;
        RECT 9.930 -0.040 10.150 0.560 ;
        RECT 10.420 0.490 12.140 0.560 ;
        RECT 10.420 0.460 11.270 0.490 ;
        RECT 10.960 0.390 11.270 0.460 ;
        RECT 11.710 0.430 12.140 0.490 ;
        RECT 13.330 0.730 13.550 1.060 ;
        RECT 13.970 0.730 14.310 0.810 ;
        RECT 14.710 0.730 15.140 0.830 ;
        RECT 13.330 0.560 15.140 0.730 ;
        RECT 13.330 0.360 13.550 0.560 ;
        RECT 13.970 0.480 14.310 0.560 ;
        RECT 14.710 0.430 15.140 0.560 ;
        RECT 16.330 0.730 16.550 1.060 ;
        RECT 17.220 1.020 17.630 1.450 ;
        RECT 19.250 1.060 19.640 1.990 ;
        RECT 22.100 1.060 22.490 1.990 ;
        RECT 22.850 1.060 23.240 1.990 ;
        RECT 24.200 1.380 24.540 1.420 ;
        RECT 25.660 1.380 26.110 1.530 ;
        RECT 24.200 1.180 26.110 1.380 ;
        RECT 24.200 1.080 24.540 1.180 ;
        RECT 25.660 1.100 26.110 1.180 ;
        RECT 26.500 1.060 26.890 1.990 ;
        RECT 27.250 1.060 27.640 1.990 ;
        RECT 33.650 1.060 34.040 1.990 ;
        RECT 17.270 1.000 17.580 1.020 ;
        RECT 16.830 0.730 17.060 0.770 ;
        RECT 16.330 0.560 17.060 0.730 ;
        RECT 16.330 0.360 16.550 0.560 ;
        RECT 16.830 0.530 17.060 0.560 ;
        RECT 17.270 0.760 17.540 1.000 ;
        RECT 17.710 0.760 18.140 0.830 ;
        RECT 17.270 0.510 18.140 0.760 ;
        RECT 17.710 0.430 18.140 0.510 ;
        RECT 19.330 0.730 19.550 1.060 ;
        RECT 19.330 0.590 20.790 0.730 ;
        RECT 22.160 0.590 22.430 1.060 ;
        RECT 19.330 0.560 22.430 0.590 ;
        RECT 19.330 0.360 19.550 0.560 ;
        RECT 20.620 0.420 22.430 0.560 ;
        RECT 13.240 0.060 13.670 0.360 ;
        RECT 16.240 0.060 16.670 0.360 ;
        RECT 19.240 0.060 19.670 0.360 ;
        RECT 9.080 -0.340 9.510 -0.040 ;
        RECT 9.840 -0.340 10.270 -0.040 ;
        RECT 21.090 -0.210 21.540 0.030 ;
        RECT 22.160 -0.040 22.430 0.420 ;
        RECT 22.930 0.730 23.150 1.060 ;
        RECT 22.930 0.560 25.260 0.730 ;
        RECT 22.930 -0.040 23.150 0.560 ;
        RECT 24.860 0.320 25.260 0.560 ;
        RECT 26.560 0.300 26.830 1.060 ;
        RECT 25.970 0.130 26.830 0.300 ;
        RECT 20.650 -0.250 21.540 -0.210 ;
        RECT 20.150 -0.380 21.540 -0.250 ;
        RECT 22.080 -0.340 22.510 -0.040 ;
        RECT 22.840 -0.340 23.270 -0.040 ;
        RECT 20.150 -0.440 20.820 -0.380 ;
        RECT 21.090 -0.400 21.540 -0.380 ;
        RECT 8.490 -0.820 8.780 -0.560 ;
        RECT 20.150 -0.600 20.530 -0.440 ;
        RECT 25.970 -0.560 26.160 0.130 ;
        RECT 26.560 -0.040 26.830 0.130 ;
        RECT 27.330 0.730 27.550 1.060 ;
        RECT 27.330 0.630 27.990 0.730 ;
        RECT 28.360 0.670 28.670 0.700 ;
        RECT 29.110 0.670 29.540 0.830 ;
        RECT 28.360 0.630 29.540 0.670 ;
        RECT 27.330 0.560 29.540 0.630 ;
        RECT 27.330 -0.040 27.550 0.560 ;
        RECT 27.820 0.490 29.540 0.560 ;
        RECT 27.820 0.460 28.670 0.490 ;
        RECT 28.360 0.390 28.670 0.460 ;
        RECT 29.110 0.430 29.540 0.490 ;
        RECT 33.730 0.730 33.950 1.060 ;
        RECT 34.230 0.740 34.460 0.770 ;
        RECT 34.230 0.730 34.640 0.740 ;
        RECT 33.730 0.560 34.640 0.730 ;
        RECT 33.730 0.360 33.950 0.560 ;
        RECT 34.230 0.530 34.460 0.560 ;
        RECT 33.640 0.060 34.070 0.360 ;
        RECT 26.480 -0.340 26.910 -0.040 ;
        RECT 27.240 -0.340 27.670 -0.040 ;
        RECT 25.890 -0.820 26.180 -0.560 ;
      LAYER met1 ;
        RECT 17.190 1.000 17.650 1.470 ;
        RECT 24.160 1.050 24.580 1.450 ;
        RECT 0.650 0.770 0.950 0.800 ;
        RECT 0.650 0.490 1.120 0.770 ;
        RECT 3.790 0.640 4.170 0.980 ;
        RECT 7.420 0.670 7.910 0.780 ;
        RECT 10.900 0.670 11.340 0.740 ;
        RECT 0.950 0.370 1.120 0.490 ;
        RECT 3.870 0.370 4.140 0.410 ;
        RECT 0.950 0.130 4.140 0.370 ;
        RECT 7.420 0.370 11.340 0.670 ;
        RECT 13.940 0.450 14.340 0.840 ;
        RECT 16.780 0.480 17.090 0.820 ;
        RECT 24.820 0.670 25.310 0.780 ;
        RECT 28.300 0.670 28.740 0.740 ;
        RECT 7.420 0.280 7.910 0.370 ;
        RECT 3.870 0.120 4.140 0.130 ;
        RECT 7.100 -0.220 7.460 0.140 ;
        RECT 16.880 -0.200 17.050 0.480 ;
        RECT 24.820 0.370 28.740 0.670 ;
        RECT 34.180 0.480 34.490 0.820 ;
        RECT 24.820 0.280 25.310 0.370 ;
        RECT 34.280 -0.200 34.450 0.480 ;
        RECT 11.010 -0.340 17.050 -0.200 ;
        RECT 8.450 -0.660 8.820 -0.530 ;
        RECT 11.010 -0.660 11.180 -0.340 ;
        RECT 20.090 -0.640 20.580 -0.220 ;
        RECT 28.410 -0.340 34.450 -0.200 ;
        RECT 8.450 -0.800 11.180 -0.660 ;
        RECT 25.850 -0.660 26.220 -0.530 ;
        RECT 28.410 -0.660 28.580 -0.340 ;
        RECT 25.850 -0.800 28.580 -0.660 ;
        RECT 8.450 -0.850 8.820 -0.800 ;
        RECT 25.850 -0.850 26.220 -0.800 ;
      LAYER met2 ;
        RECT 17.190 1.340 17.650 1.470 ;
        RECT 14.010 1.070 17.650 1.340 ;
        RECT 3.790 0.690 4.170 0.980 ;
        RECT 14.010 0.840 14.270 1.070 ;
        RECT 17.190 1.000 17.650 1.070 ;
        RECT 24.160 1.050 24.580 1.450 ;
        RECT 3.790 0.640 7.100 0.690 ;
        RECT 4.020 0.550 7.100 0.640 ;
        RECT 6.950 0.140 7.100 0.550 ;
        RECT 13.940 0.450 14.340 0.840 ;
        RECT 6.950 -0.220 7.460 0.140 ;
        RECT 7.210 -0.810 7.410 -0.220 ;
        RECT 20.090 -0.640 20.580 -0.220 ;
        RECT 20.240 -0.810 20.410 -0.640 ;
        RECT 24.160 -0.810 24.360 1.050 ;
        RECT 7.210 -0.950 24.360 -0.810 ;
  END
END dff
END LIBRARY

