* Assignment 1, Q2: INVX2 CMOS Inverter - Transient Analysis

.lib ~/VLSI_Design/open_pdks/sources/sky130_fd_pr/models/sky130.lib.spice tt

* parameters
.param VDD=1.8
.param Lmin=0.15
.param Wn1=0.42
.param Wp1=1.31   ; INVX1 widths
.param Wn2=0.84
.param Wp2=2.62   ; INVX2 widths = 2 * INVX1

.param ASn1=Wn1*0.3
.param ADn1=Wn1*0.3
.param PSn1=2*(Wn1+0.3)
.param PDn1=2*(Wn1+0.3)

.param ASp1=Wp1*0.3
.param ADp1=Wp1*0.3
.param PSp1=2*(Wp1+0.3)
.param PDp1=2*(Wp1+0.3)

.param ASn2=Wn2*0.3
.param ADn2=Wn2*0.3
.param PSn2=2*(Wn2+0.3)
.param PDn2=2*(Wn2+0.3)

.param ASp2=Wp2*0.3
.param ADp2=Wp2*0.3
.param PSp2=2*(Wp2+0.3)
.param PDp2=2*(Wp2+0.3)

Vdd vdd gnd DC {VDD}
Vin in gnd PULSE(0 {VDD} 0p 20p 20p 1n 2n)

* Main Circuit
Xinv2 in vdd gnd out INVX2_sub
Xload out vdd gnd out_load INVX1_sub

* Sub - Ckt Defn
.subckt INVX1_sub a vdd vss z
* NMOS
XM1 z a vss vss sky130_fd_pr__nfet_01v8 L={Lmin} W={Wn1} AS={ASn1} AD={ADn1} PS={PSn1} PD={PDn1}
* PMOS
XM2 z a vdd vdd sky130_fd_pr__pfet_01v8 L={Lmin} W={Wp1} AS={ASp1} AD={ADp1} PS={PSp1} PD={PDp1}
.ends INVX1_sub

.subckt INVX2_sub a vdd vss z
* NMOS
XM1 z a vss vss sky130_fd_pr__nfet_01v8 L={Lmin} W={Wn2} AS={ASn2} AD={ADn2} PS={PSn2} PD={PDn2}
* PMOS
XM2 z a vdd vdd sky130_fd_pr__pfet_01v8 L={Lmin} W={Wp2} AS={ASp2} AD={ADp2} PS={PSp2} PD={PDp2}
.ends INVX2_sub


.tran 1ps 10ns 0 10p
.param Vhalf={VDD/2}
.meas tran tr TRIG v(out) VAL='0.1*VDD' RISE=1 TARG v(out) VAL='0.9*VDD' RISE=1
.meas tran tf TRIG v(out) VAL='0.9*VDD' FALL=1 TARG v(out) VAL='0.1*VDD' FALL=1
.meas tran tpHL TRIG v(in) VAL='Vhalf' RISE=1 TARG v(out) VAL='Vhalf' FALL=1
.meas tran tpLH TRIG v(in) VAL='Vhalf' FALL=1 TARG v(out) VAL='Vhalf' RISE=1

.control
run
print tran tr tf tpHL tpLH
print param Wn2 Wp2
plot v(in) v(out)
.endc

.end

